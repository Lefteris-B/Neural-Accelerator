module wishbone_slave
(
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,  // Assuming 4-bit select lines for Wishbone
    input [31:0] wbs_dat_i, // Assuming 32-bit data width for Wishbone
    input [31:0] wbs_adr_i, // Assuming 32-bit address width for Wishbone
    output reg wbs_ack_o,
    output reg [31:0] wbs_dat_o, // Data to be read by the master
    output reg wbs_rdy_o
);

    // Parameters
    parameter Rows = 8; // Placeholder value
    parameter Columns = 8; // Placeholder value
    parameter Width = 8; // 8-bit signed numbers
    parameter AddressRange = 32; // Placeholder value. This defines how many registers or memory locations the slave has.

    // Internal Registers (Assuming 32-bit registers for simplicity. Adjust size accordingly.)
    reg [31:0] internal_registers[AddressRange-1:0];
    reg [31:0] temp_data;

    // Control FSM states
    typedef enum {
        IDLE,
        READ,
        WRITE
    } fsm_state_t;

    fsm_state_t current_state, next_state;

    // Control FSM
    always @(posedge wb_clk_i or negedge wb_rst_i) begin
        if (!wb_rst_i) begin
            current_state <= IDLE;
        end else begin
            current_state <= next_state;
        end
    end

    // FSM Logic
    always @(current_state or wbs_stb_i or wbs_cyc_i or wbs_we_i or wbs_adr_i or wbs_dat_i) begin
        case (current_state)
            IDLE: begin
                wbs_ack_o = 0;
                if (wbs_stb_i && wbs_cyc_i) begin
                    if (wbs_we_i) begin
                        temp_data = wbs_dat_i;
                        next_state = WRITE;
                    end else begin
                        wbs_dat_o = internal_registers[wbs_adr_i];
                        next_state = READ;
                    end
                end else begin
                    next_state = IDLE;
                end
            end

            READ: begin
                wbs_ack_o = 1;
                wbs_rdy_o = 1; // Ready to accept new requests
                next_state = IDLE;
            end

            WRITE: begin
                internal_registers[wbs_adr_i] = temp_data;
                wbs_ack_o = 1;
                wbs_rdy_o = 1; // Ready to accept new requests
                next_state = IDLE;
            end

            default: begin
                wbs_ack_o = 0;
                wbs_rdy_o = 0;
                next_state = IDLE;
            end
        endcase
    end

endmodule
